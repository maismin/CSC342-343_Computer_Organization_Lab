-- library declaration
library IEEE;
use IEEE.std_logic_1164.all;

-- entity
entity test_4b_fadder is
end test_4b_fadder;

-- architecture
architecture arch_test of test_4b_fadder is
  -- component
  -- 4 bit full adder ---------------------------
  component mai_four_bit_full_adder
  port (  X, Y : in std_logic_vector(3 downto 0);
          Cin  : in std_logic;
          Sum  : out std_logic_vector(3 downto 0);
          Cout : out std_logic);
  end component;

  -- intermediate signal declarations
  signal t_x, t_y, t_sum  : std_logic_vector(3 downto 0);
  signal t_cin, t_cout    : std_logic;
  signal error            : std_logic := '0';
  
begin
  t:  mai_four_bit_full_adder port map(X => t_x, Y => t_y, Cin => t_cin, Sum => t_sum, Cout => t_cout);
  process
  begin
    t_cin <= '0';
    t_x <= "0000";
    t_y <= "0000";
    wait for 1 ns;
    if (t_sum /= "0000" or t_cout /= '0') then
      error <= '1';
    end if;
    
    wait for 200 ns;
    t_cin <= '1';
    t_x <= "1111";
    t_y <= "1111";
    wait for 1 ns;
    if (t_sum /= "1111" or t_cout /= '1') then
      error <= '1';
    end if;
    
    wait for 200 ns;
    t_cin <= '0';
    t_x <= "1111";
    t_y <= "1111";
    wait for 1 ns;
    if (t_sum /= "1110" or t_cout /= '1') then
      error <= '1';
    end if;
    
    wait for 200 ns;
    t_cin <= '1';
    t_x <= "1111";
    t_y <= "0111";
    wait for 1 ns;
    if (t_sum /= "0111" or t_cout /= '1') then
      error <= '1';
    end if;
    
    wait for 200 ns;
    t_cin <= '1';
    t_x <= "1010";
    t_y <= "0101";
    wait for 1 ns;
    if (t_sum /= "0000" or t_cout /= '1') then
      error <= '1';
    end if;
    
    wait for 200 ns;
    t_cin <= '1';
    t_x <= "1001";
    t_y <= "0000";
    wait for 1 ns;
    if (t_sum /= "1010" or t_cout /= '0') then
      error <= '1';
    end if;
    
    wait for 200 ns;
    t_cin <= '1';
    t_x <= "1100";
    t_y <= "0011";
    wait for 1 ns;
    if (t_sum /= "0000" or t_cout /= '1') then
      error <= '1';
    end if;
    
    wait for 200 ns;
      
    if (error = '0') then
      report "No errors detected. Simulation successful" severity failure;
    else
      report "Error detected" severity failure;
    end if;
  end process;
end arch_test;
